66
34
0
